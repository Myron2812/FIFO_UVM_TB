`define DATA_W 128
